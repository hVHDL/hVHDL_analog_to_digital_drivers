library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package sigma_delta_cic_filter_pkg is

end package sigma_delta_cic_filter_pkg;

package body sigma_delta_cic_filter_pkg is

end package body sigma_delta_cic_filter_pkg;
